module instruction_memory (
    
);
    // .a(instr_mem_if.pc[11:2]),
    // .spo(instr_mem_if.instr)

endmodule