`timescale 1ns/1ps

module mem_wb_reg (

);
    
endmodule