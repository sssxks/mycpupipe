`timescale 1ns/1ps
`default_nettype none

module instruction_memory_impl (
    input wire [9:0] a,
    output wire [31:0] spo
);
    
endmodule