`timescale 1ns/1ps

module id_ex_reg (
    logic clk,
    logic reset,

    
);
    
endmodule