`timescale 1ns/1ps
`default_nettype none

module data_memory_impl(
    input wire clka,
    input wire [3:0] wea,
    input wire [9:0] addra,
    input wire [31:0] dina,
    output wire [31:0] douta
);
    
endmodule