
// typedef struct {
    
// } id_ex_flow_t;