`timescale 1ns/1ps

module id_ex_reg (
    input logic clk,
    input logic reset
);
    
endmodule