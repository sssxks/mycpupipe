module my_data_memory (
    input logic clk,
    data_memory_if.mem mem_if
);
    
endmodule