module my_data_memory (
    
);
    
endmodule