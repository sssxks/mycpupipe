`timescale 1ns/1ps

module ex_mem_reg (
);
    
endmodule